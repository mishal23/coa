//Mishal Shah
//16CO125
//Random message generation
//16 Oct 2017

module A(output reg[3:0] message_out,input[3:0][3:0] message_in,input clock);
    reg[3:0] rnd=3'b000;                         //random is set as 0
    always@(posedge clock) begin
        if(rnd==3'b000) begin
            rnd <= {$random}%16+1;               //random is changed
            message_out <= {$random}%8;          //random msg sent by A
            $display("Time:%0t\nA sent %b to B",$time,message_out);         //msg displayed
            $display("B responded with %b %b %b %b\n",message_in[0],message_in[1],message_in[2],message_in[3]);    //msg recieved displayed                            
        end 
        else begin
            rnd <= rnd - 1;  //random variable decremented to send msg at random interval
        end
        
    end
endmodule

module B(output reg[3:0][3:0] message_out,input[3:0] message_in,input clock);
    always@(posedge clock) begin
        if(message_in !== 4'bzzzz) begin
            message_out[0] <= {$random}%16;            //random msg generated by B
            message_out[1] <= {$random}%16;
            message_out[2] <= {$random}%16;
            message_out[3] <= {$random}%16;
        end
    end
endmodule